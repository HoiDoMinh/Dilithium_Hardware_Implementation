`timescale 1ns/1ps

module tb_polyvec_matrix_pointwise_montgomery;

  reg clock;
  reg reset;
  reg start;

  reg  signed [40959:0] v_in;    // polyvecl v (5 ?a th?c, m?i 8192b)
  reg  signed [65535:0] mat1;    // d? li?u ma tr?n n�n
  reg  signed [65535:0] mat2;
  reg  signed [65535:0] mat3;
  reg  signed [49151:0] mat4;

  wire signed [49151:0] t_out;   // 6 ?a th?c k?t qu? (6�8192b)
  wire done;

  integer i, j;

  polyvec_matrix_pointwise_montgomery dut (
      .clock(clock),
      .reset(reset),
      .start(start),
      .v_in(v_in),
      .mat1(mat1),
      .mat2(mat2),
      .mat3(mat3),
      .mat4(mat4),
      .t_out(t_out),
      .done(done)
  );


  initial clock = 0;
  always #5 clock = ~clock;


  initial begin
    reset = 1;
    start = 0;
    v_in  = 0;
    mat1  = 0;mat2  = 0;mat3  = 0;mat4  = 0;

    #20 reset = 0;

    for (i = 0; i < 256; i = i + 1) begin

      v_in[(i*32) +: 32] = i + 1;
    end
/*
    for (i = 0; i < 2048; i = i + 1) begin
      mat1[(i*32) +: 32] = 1000 + i;   // ch? c?n gi� tr? m?u
      mat2[(i*32) +: 32] = 2000 + i;
      mat3[(i*32) +: 32] = 3000 + i;
    end
    for (i = 0; i < 1536; i = i + 1) begin
      mat4[(i*32) +: 32] = 4000 + i;
    end
*/

    #10 start = 1;

    wait(done == 1);
    #10 start = 0;

    for (i = 0; i < 6; i = i + 1) begin
      $display("---- t[%0d] ----", i);
      for (j = 0; j < 8; j = j + 1) begin
        // ch? in 8 h? s? ??u m?i ?a th?c cho ng?n
        $display("  coeff[%0d] = %d",
                 j, $signed(t_out[8192*i + (j*32) +: 32]));
      end
    end

    #50 $finish;
  end

endmodule

