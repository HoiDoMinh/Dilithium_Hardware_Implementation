`timescale 1ns/1ps
`include "byte_and_print.vh"

module tb_pack_pk;
    reg  [255:0]      rho_in;
    reg  [49151:0]    t1_in;
    wire [15615:0]    pk_out;

    pack_pk dut(
        .rho_in(rho_in),
        .t1_in(t1_in),
        .pk_out(pk_out)
    );


    wire [7:0] pk_bytes [0:1951];

    integer i;

    `BYTE_ASSIGN_GEN(PKMAP, 1952, pk_out, pk_bytes)


    initial begin

        // RHO from C
        rho_in = 256'h449e6340f762807b7675c26c548f69d84e7c623176dc341ee7bc8bc4b13f77e5;

        // T1 from C (49152 bits)
        t1_in  = 49152'h000003a20000035600000069000003ce000000b3000003e90000035f000000840000036900000345000003f2000001400000004d000003ef00000389000003c20000035b00000290000003ab000001b50000037b00000023000001890000010e000002fe0000022b000002dd00000083000003a4000003970000026700000200000001470000034000000103000003b2000000dd0000024e00000296000001dc000002b90000011000000035000001340000007300000042000003460000001600000142000001e60000009d000000440000003200000302000003b80000028a000000a1000000a8000002340000004400000377000002e10000003800000280000002e9000002e4000003c10000035d00000113000000d0000002bc0000000e000000e5000001b20000037e000003be00000089000003bf000000b0000003d70000010d000002b50000039a000000fe000003bc00000385000000c5000002e2000001c5000003e500000299000001340000037e000001180000030f0000002400000202000001790000030f0000010a000003d6000001a40000016200000266000002d30000028c000002d2000003e4000003ce00000276000003db000002db000002f0000000940000025a000001a20000020600000348000003ab0000034d000002290000022a0000017e000003e1000003940000022b000002ab000003b500000362000003fa000000fe0000024f0000033a00000198000002140000006600000012000000ae00000146000001d7000003d50000001e0000009e000001c2000001c5000003df00000112000002fc0000026c000002a9000002c600000096000003ec000000d6000000b10000002c000001d50000006a000001280000034500000025000001db00000295000002ed0000021f000002ba000000d20000025300000269000002a6000000ec0000024f000000780000032b00000363000003ee0000021a000000d300000271000001750000008e000000f500000399000001cf000001f6000001b50000013e00000067000002f800000374000003f200000009000003ac000002470000027f00000032000000c10000026b00000210000000c7000001be000002440000006b0000028200000268000002e5000000c6000000dd000003060000032b0000009a0000012a000003f20000027600000155000003c2000002b800000208000000d700000383000001f7000000a9000003b6000001b500000261000000620000005e0000020400000114000002d6000000420000034f000001e00000036c00000139000001350000015f0000026b000001e6000000d60000039700000291000001ee0000038c00000267000003ce0000032f0000035e0000028c0000039e0000038e0000019b000003fe00000070000000160000000b000001d4000003620000014d0000014f00000260000003ca000003040000036d000003cf0000006e000002d8000003ef0000022f000000bf0000010b0000025e000002140000029d0000007f000002eb000000f40000015d0000026d0000033a0000023200000270000003d80000017800000191000001eb00000280000003e3000001e80000016f000002ff0000033c000000db0000020d000003e4000001d6000002450000010f0000016a00000134000001b8000000cd000003ef000003f6000003ac0000031a000000ac00000001000000ea00000168000002bb0000022b00000117000002c10000018c000001f10000032e000002f300000227000003100000033800000289000001a9000001bb00000148000001c900000182000001e70000023a000000db000000c400000369000003f4000000da00000099000000f30000000100000044000000f5000003240000023500000193000003d400000389000000900000024200000394000001190000005e00000373000001820000002a00000112000001410000027700000347000000760000032f0000019b000002ca000000f700000133000000bc000001b10000013e00000354000000e3000003fd000000a7000001b7000002320000029d00000352000001ac0000011d0000029600000217000002a5000002e0000003f700000190000002b500000245000003a5000002f8000001fa00000042000002d9000003f5000002af000001850000024b0000031300000240000002a40000035b0000020a000002360000019e000000db000000870000036400000050000001eb000003d100000083000001cc000000f3000001cb000002c900000106000003f300000302000001620000017b000002e10000002f0000028400000265000001890000002a000001ca000001390000024a000002bc0000035500000207000003c6000003600000030e000001ab00000052000003e70000036000000095000000ab000003b5000002c3000001bc0000018700000361000001d00000001d000001cf000001e7000003d600000059000003c800000170000001e0000001bd0000004100000074000002f30000017c0000022c000003090000007200000355000001f50000014d000003af000001ae0000016b000001ad00000068000001bf00000290000000e8000000340000021b00000205000001cd000001730000003000000278000002a700000208000001160000028f00000084000003840000034f000001ea00000158000001b6000000a9000000330000032d0000000e000003c1000000c4000000da0000033e0000008200000056000001600000012900000085000000d300000384000003c20000036f0000008500000202000001a00000038d0000032f000001c600000196000003d200000365000001d2000001ef0000020b000003da00000014000000980000013e000003cb000003260000011d0000035900000214000000ce00000034000003e10000000200000220000003ce00000021000003e40000035a000001b2000000a20000030d0000017c00000397000003cb000001ba0000037b0000022e000002bb000003360000038d0000002b00000214000000ed000003c80000027a00000322000002420000022d000002b400000184000003c4000000310000036c000003ef00000384000003f3000003600000026f00000254000002c5000001d00000015f000000a600000302000002f2000002190000033b000002c1000002ec0000037900000276000002ff0000031b0000011400000242000000db000002310000010f0000039d000000b1000001e2000002d1000003eb000001680000009a0000017700000361000003410000021d000000600000039c0000039b0000037d0000034f000000d5000003cc00000093000000ba000003c50000019f0000024a000002ae0000031d000000bc00000372000002ce000001bb0000007e000002dd0000014c000003a6000003630000032800000179000000ae0000031a00000092000003f5000003f6000001a90000008400000065000002ff0000002400000209000001b400000370000002cd000000df0000012d000003f1000003bb0000007d0000007100000285000002de000002ec00000052000002cf000002ec000002d6000001d800000080000001ac000001ce000001a3000003eb000002e9000002bc0000026e000000b600000222000003a7000000cf00000146000003a80000020d0000023300000309000001880000017600000233000002390000019c00000235000003dd000000e7000002b40000021c00000142000003bc0000021000000020000002e400000394000000a200000298000002000000011300000231000003640000027f000002100000028000000173000001db0000011500000228000000d50000013400000109000002f90000020b00000215000001f3000003f9000001ef000001990000006a000003740000009b000000cb00000220000003010000029b000003b10000025d00000328000000c6000000050000004f0000035a0000034a000003660000008d000002df00000341000003b8000000c2000003bb000000f60000032400000301000001f60000028d000000ed000001190000028b0000032b00000346000003b5000000970000018e000001c0000001b50000035a000003f7000003900000035000000281000000390000026a000000c80000029f000001c70000008f000001c1000001100000029b00000294000003a80000030c000003f2000001a3000003fe000003e0000003a500000243000000b3000000a00000003c000002050000001600000155000000fd000002ad00000241000003070000028a00000298000001360000029d000001d8000001c1000000c600000190000001a90000001a000000b90000025300000360000001710000027200000159000002770000012900000171000000a8000003dc000001180000031a000003940000020700000260000001db0000029e000002af0000005b0000031c000001330000021c0000014a000000e70000038600000018000001b7000002be00000281000001ea000001090000018500000361000002d1000003fb0000028b00000213000003830000034a0000036f0000005e0000003900000343000002870000022f000001da000001cf000003f70000026300000307000000b7000001e10000022a0000014400000321000000f90000009600000086000002a800000204000002fc00000299000003a00000002e000003e500000313000003070000034d000001ac000002aa000001080000014f000000940000019500000146000001d9000001ea00000360000001e3000003030000038e0000021a0000018c0000027e000000a90000019d0000013700000385000002240000023d000002f400000054000002f40000009d000003e4000003650000017f0000003b0000027f000001da00000133000001cb000001d000000398000001f8000001750000016b00000166000000ba00000167000000ce000003b600000360000002b500000082000001ac0000022c0000036d0000009e000000390000027b0000020000000097000000f000000282000001da0000008500000117000002a0000001500000010d000001d0000000a40000019d00000293000003f4000000b2000003030000035d000001f000000361000003000000016b000002bf0000001b0000009b000001e1000003630000036600000068000000b8000003f300000258000001fb0000027c000000130000018f0000021c000003f0000001bf0000003e000001d300000014000003e600000334000003c800000165000002060000014800000231000002d9000002c30000034e0000038b000001b700000294000002cf000003a7000000b7000003f9000000d5000002920000029b00000118000003d400000200000001ba00000104000000230000013a00000003000003370000015500000011000000c800000003000001a5000003bd0000032d0000033400000360000001c00000019d00000233000000a5000000a6000003e200000176000001470000001b000000d9000001ce000000fd0000030100000303000002ac000002a400000218000001320000014e00000215000003600000028100000151000000030000025100000257000001d300000351000000740000013d0000035200000023000002fb000001c90000032f000001d70000011e000002960000026a000002e10000008d00000298000000e50000037f0000002b000000fc000001730000031e0000023f00000278000001010000002f000003430000006d0000036a000000ee000000e9000000660000030d0000028400000324000003b00000032c000001e60000001b000002fa000003f5000003d900000350000001d4000002c70000016f000000d30000008a00000028000000510000025e000002c50000032a0000020a000001a90000015a0000011e000002b10000030200000115000000b9000001c8000002f00000007200000053000003450000010d0000037c0000019a000002830000028900000213000000af0000009c0000017a00000262000000000000033e0000019e000002460000002a0000019f0000002e00000088000001fc000000d2000000660000010400000176000003a300000340000001b7000000c80000003f0000019d000000a0000002170000002c0000032d0000038e00000049000002ff000000cd0000008b0000035600000236000002c0000001150000023a0000009100000232000001e8000001100000003c0000016800000251000001c90000004c00000149000002670000009b000002370000012a000003f8000002440000022d0000003f00000070000000da000001c1000003ad00000252000003ac000001990000034b000002b9000001050000025a000003950000004100000226000003ca0000001c0000000d0000025b00000122000003a400000062000003e10000003f0000023f000001310000033c0000024b0000017a0000015100000180000001ab00000037000001680000014a0000020a00000341000001f8000002cb0000017b00000188000000a7000003ea000000140000006e00000367000003ad000001b40000021e0000024c00000214000001d1000003640000012600000150000000a8000000c6000002e30000000100000178000003e20000026800000272000002b3000003c1000000f700000303000003b200000187000001a00000028700000050000001120000031e00000385000001170000035e0000007e000002a4000000890000002e0000024b000001af0000034d000003b3000000e80000035e000000dc000002210000023800000315000000970000037c00000132000002ac0000038c000003f2000002bb000001060000031200000264000002c0000002560000002b000001c40000002700000031000000450000032f00000312000002b000000313000000a600000308000000b70000035f0000016d0000002a000001dc000003050000026a00000310000000c90000015900000133000003470000014600000143000003b6000003f400000240000001600000022500000392000002a90000003600000246000001820000022b0000037e0000009e000002e000000288000002fe0000003300000287000002b50000005800000016000000d700000136000003fa00000150000000d200000237000003b50000000c0000022a0000003e00000158000003240000002e0000014e00000093000000d1000000910000006400000004000000b00000002e00000269000000d7000002700000030b000002d4000003b3000002a3000003a200000185000000b000000060000001ce0000019d000002960000035b0000009e000002b2000003b60000011300000321000003410000018b000003dd000003b700000238000002f2000002270000008500000116000002e2000000c3000003d40000038e0000013f000002430000037700000238000001a400000077000001340000031300000172000001bb0000007a0000020500000274000001a7000002f80000034000000045000002c7000001c3000001120000017a00000282000003c50000011f0000020b000003eb0000023800000354000001a2000001cf000002f3000002b30000016b00000301000002bc000003620000004d0000010d0000014500000174000001e5000003c5000002350000008c0000037000000187000003f700000266000003f600000180000002dc0000005a0000026e0000034d00000249000002f40000005d000001940000011a0000029c000002a1000002a0000000e50000028c000000dd0000015e0000003100000233000001f4000000850000014400000009000001dc0000030a000002d10000015c0000012c0000000f000000bd000002e4000000f50000015e00000001000001a7000003a8000000bb000001f800000036000001280000030c0000001e00000238000003440000019b0000033d0000034b000000e0000003b9000000d80000030b00000383000001b40000000e0000023d000002e30000002c000002f800000194000002de00000289000001cb0000022c000001d80000006500000124000001470000019d000000960000016d000000a3000001590000032a00000340000001ea000003e9000002a9000003810000011700000270000000180000002d00000104000002a1000000e6000003fc000001a200000039000000a300000106000002d200000193000000690000000a000002ec00000332000002b000000143000000f60000014f000002c8000000870000019200000015000002190000027600000378000003b4000001be000000e10000014100000179000001c30000026e000003d40000029f000000a8000002a0000000ed000002150000008e0000020700000160000001d300000213000003ec0000025800000036000002500000026c000000bb000003e90000009000000140000000470000029600000089000001d500000162000002620000035400000319000003400000009c000000da000003da00000017;


        #10;

        `PRINT_HEX_ARRAY("pk_out (Verilog)", pk_bytes, 1952)

        $finish;
    end

endmodule
