
//a=a1?*2^D+a0?                 D=13    

module power2round(
    input signed [31:0] a,
    output signed [31:0] a0,
    output signed [31:0] a1
);
    localparam D = 13;
    
    assign a1 = (a + (1 << (D-1))-1) >>> D;  // Signed shift
    assign a0 = a - (a1 << D);
    
endmodule
