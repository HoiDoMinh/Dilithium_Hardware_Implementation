`timescale 1ns/1ps
`include "byte_and_print.vh"

module tb_polyz_pack;

  // a_in n�n l� wire n?u d�ng assign
  wire [8191:0] a_in;
  wire [5119:0] r_out;
  integer i;
  assign a_in = 8192'hffffb34d00007a0affffb3e700007914ffffb4810000781effffb51b00007728ffffb5b500007632ffffb64f0000753cffffb6e900007446ffffb78300007350ffffb81d0000725affffb8b700007164ffffb9510000706effffb9eb00006f78ffffba8500006e82ffffbb1f00006d8cffffbbb900006c96ffffbc5300006ba0ffffbced00006aaaffffbd87000069b4ffffbe21000068beffffbebb000067c8ffffbf55000066d2ffffbfef000065dcffffc089000064e6ffffc123000063f0ffffc1bd000062faffffc25700006204ffffc2f10000610effffc38b00006018ffffc42500005f22ffffc4bf00005e2cffffc55900005d36ffffc5f300005c40ffffc68d00005b4affffc72700005a54ffffc7c10000595effffc85b00005868ffffc8f500005772ffffc98f0000567cffffca2900005586ffffcac300005490ffffcb5d0000539affffcbf7000052a4ffffcc91000051aeffffcd2b000050b8ffffcdc500004fc2ffffce5f00004eccffffcef900004dd6ffffcf9300004ce0ffffd02d00004beaffffd0c700004af4ffffd161000049feffffd1fb00004908ffffd29500004812ffffd32f0000471cffffd3c900004626ffffd46300004530ffffd4fd0000443affffd59700004344ffffd6310000424effffd6cb00004158ffffd76500004062ffffd7ff00003f6cffffd89900003e76ffffd93300003d80ffffd9cd00003c8affffda6700003b94ffffdb0100003a9effffdb9b000039a8ffffdc35000038b2ffffdccf000037bcffffdd69000036c6ffffde03000035d0ffffde9d000034daffffdf37000033e4ffffdfd1000032eeffffe06b000031f8ffffe10500003102ffffe19f0000300cffffe23900002f16ffffe2d300002e20ffffe36d00002d2affffe40700002c34ffffe4a100002b3effffe53b00002a48ffffe5d500002952ffffe66f0000285cffffe70900002766ffffe7a300002670ffffe83d0000257affffe8d700002484ffffe9710000238effffea0b00002298ffffeaa5000021a2ffffeb3f000020acffffebd900001fb6ffffec7300001ec0ffffed0d00001dcaffffeda700001cd4ffffee4100001bdeffffeedb00001ae8ffffef75000019f2fffff00f000018fcfffff0a900001806fffff14300001710fffff1dd0000161afffff27700001524fffff3110000142efffff3ab00001338fffff44500001242fffff4df0000114cfffff57900001056fffff61300000f60fffff6ad00000e6afffff74700000d74fffff7e100000c7efffff87b00000b88fffff91500000a92fffff9af0000099cfffffa49000008a6fffffae3000007b0fffffb7d000006bafffffc17000005c4fffffcb1000004cefffffd4b000003d8fffffde5000002e2fffffe7f000001ecffffff19000000f6ffffffb300000000;

  polyz_pack dut (
    .a_in(a_in),
    .r_out(r_out)
  );

  wire [7:0] r_out_t [0:639];
  `BYTE_ASSIGN_GEN(r, 640, r_out, r_out_t)

  initial begin
    #1;
    `PRINT_HEX_ARRAY("r out", r_out_t, 640)
    $finish;
  end

endmodule

