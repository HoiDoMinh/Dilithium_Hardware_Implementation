`timescale 1ns/1ps

module tb_randombytes;
    parameter in_len = 32;
    reg clk, rst_n, start;
    wire [in_len*8-1:0] zeta_out;
    wire random_done;

    randombytes #(.IN_LEN(in_len)) uut (
        .clk(clk),
        .rst_n(rst_n),
        .start(start),
        .zeta_out(zeta_out),
        .random_done(random_done)
    );

    // clock 10 ns period
    always #5 clk = ~clk;

    initial begin
        clk = 0;rst_n = 0;start = 0;

        #20 rst_n = 1;         
        #10 @(posedge clk);     


        start = 1;
        @(posedge clk);
        start = 0;
        fork
            begin
                wait(random_done);
                $display("Random output = %h", zeta_out);
                #100 $finish;
            end
            begin
                #1000;
                if (!random_done) begin
                    $display("ERROR: timeout waiting for random_done");
                    $finish;
                end
            end
        join
    end
endmodule
