`timescale 1ns / 1ps

module parallel_invntt_tomont_32bit
(
    input clock,
    input reset,
    input start,
    input signed [0:8191] inp,
    output rd_ready,
    output rd_done,
    output done,
    output wr_done,
    output signed [0:8191] out
);
    localparam SIZE = 4;
    localparam IDLE = 4'd0, PRE_RD_INP = 4'd1 ,RD_INP = 4'd2, CALC_1 = 4'd3, CALC_2 = 4'd4,
               CALC_3 = 4'd5, CALC_4 = 4'd6, WR_OUT = 4'd7, DONE = 4'd8;

    reg [SIZE-1:0] state;
    reg [SIZE-1:0] next_state;

    reg signed [0:8191] temp_inp;
    reg temp_rd_ready;
    reg temp_rd_done;
    reg temp_done;
    reg temp_wr_done;
    reg signed [0:8191] temp_out;

    reg new_fqmul_32bit_start;
    wire [0:127] new_fqmul_32bit_done;
    wire new_fqmul_32bit_final_done;

    reg signed [0:4095] temp_i1;
    reg signed [0:4095] temp_i2;
    wire signed [0:4095] temp_o1;
    reg signed [0:4095] temp_o2;

    reg signed [31:0] f = 32'd41978;
    reg [8:0] len;
    reg [1:0] counter;

    integer n;
    integer m;

    reg signed [0:8191] zetas =
    {
    32'sd0, 32'sd25847, -32'sd2608894, -32'sd518909, 32'sd237124, -32'sd777960, -32'sd876248, 32'sd466468, 
    32'sd1826347, 32'sd2353451, -32'sd359251, -32'sd2091905, 32'sd3119733, -32'sd2884855, 32'sd3111497, 32'sd2680103, 
    32'sd2725464, 32'sd1024112, -32'sd1079900, 32'sd3585928, -32'sd549488, -32'sd1119584, 32'sd2619752, -32'sd2108549, 
    -32'sd2118186, -32'sd3859737, -32'sd1399561, -32'sd3277672, 32'sd1757237, -32'sd19422, 32'sd4010497, 32'sd280005, 
    32'sd2706023, 32'sd95776, 32'sd3077325, 32'sd3530437, -32'sd1661693, -32'sd3592148, -32'sd2537516, 32'sd3915439, 
    -32'sd3861115, -32'sd3043716, 32'sd3574422, -32'sd2867647, 32'sd3539968, -32'sd300467, 32'sd2348700, -32'sd539299, 
    -32'sd1699267, -32'sd1643818, 32'sd3505694, -32'sd3821735, 32'sd3507263, -32'sd2140649, -32'sd1600420, 32'sd3699596, 
    32'sd811944, 32'sd531354, 32'sd954230, 32'sd3881043, 32'sd3900724, -32'sd2556880, 32'sd2071892, -32'sd2797779, 
    -32'sd3930395, -32'sd1528703, -32'sd3677745, -32'sd3041255, -32'sd1452451, 32'sd3475950, 32'sd2176455, -32'sd1585221, 
    -32'sd1257611, 32'sd1939314, -32'sd4083598, -32'sd1000202, -32'sd3190144, -32'sd3157330, -32'sd3632928, 32'sd126922, 
    32'sd3412210, -32'sd983419, 32'sd2147896, 32'sd2715295, -32'sd2967645, -32'sd3693493, -32'sd411027, -32'sd2477047, 
    -32'sd671102, -32'sd1228525, -32'sd22981, -32'sd1308169, -32'sd381987, 32'sd1349076, 32'sd1852771, -32'sd1430430, 
    -32'sd3343383, 32'sd264944, 32'sd508951, 32'sd3097992, 32'sd44288, -32'sd1100098, 32'sd904516, 32'sd3958618, 
    -32'sd3724342, -32'sd8578, 32'sd1653064, -32'sd3249728, 32'sd2389356, -32'sd210977, 32'sd759969, -32'sd1316856, 
    32'sd189548, -32'sd3553272, 32'sd3159746, -32'sd1851402, -32'sd2409325, -32'sd177440, 32'sd1315589, 32'sd1341330, 
    32'sd1285669, -32'sd1584928, -32'sd812732, -32'sd1439742, -32'sd3019102, -32'sd3881060, -32'sd3628969, 32'sd3839961, 
    32'sd2091667, 32'sd3407706, 32'sd2316500, 32'sd3817976, -32'sd3342478, 32'sd2244091, -32'sd2446433, -32'sd3562462, 
    32'sd266997, 32'sd2434439, -32'sd1235728, 32'sd3513181, -32'sd3520352, -32'sd3759364, -32'sd1197226, -32'sd3193378, 
    32'sd900702, 32'sd1859098, 32'sd909542, 32'sd819034, 32'sd495491, -32'sd1613174, -32'sd43260, -32'sd522500, 
    -32'sd655327, -32'sd3122442, 32'sd2031748, 32'sd3207046, -32'sd3556995, -32'sd525098, -32'sd768622, -32'sd3595838, 
    32'sd342297, 32'sd286988, -32'sd2437823, 32'sd4108315, 32'sd3437287, -32'sd3342277, 32'sd1735879, 32'sd203044, 
    32'sd2842341, 32'sd2691481, -32'sd2590150, 32'sd1265009, 32'sd4055324, 32'sd1247620, 32'sd2486353, 32'sd1595974, 
    -32'sd3767016, 32'sd1250494, 32'sd2635921, -32'sd3548272, -32'sd2994039, 32'sd1869119, 32'sd1903435, -32'sd1050970, 
    -32'sd1333058, 32'sd1237275, -32'sd3318210, -32'sd1430225, -32'sd451100, 32'sd1312455, 32'sd3306115, -32'sd1962642, 
    -32'sd1279661, 32'sd1917081, -32'sd2546312, -32'sd1374803, 32'sd1500165, 32'sd777191, 32'sd2235880, 32'sd3406031, 
    -32'sd542412, -32'sd2831860, -32'sd1671176, -32'sd1846953, -32'sd2584293, -32'sd3724270, 32'sd594136, -32'sd3776993, 
    -32'sd2013608, 32'sd2432395, 32'sd2454455, -32'sd164721, 32'sd1957272, 32'sd3369112, 32'sd185531, -32'sd1207385, 
    -32'sd3183426, 32'sd162844, 32'sd1616392, 32'sd3014001, 32'sd810149, 32'sd1652634, -32'sd3694233, -32'sd1799107, 
    -32'sd3038916, 32'sd3523897, 32'sd3866901, 32'sd269760, 32'sd2213111, -32'sd975884, 32'sd1717735, 32'sd472078, 
    -32'sd426683, 32'sd1723600, -32'sd1803090, 32'sd1910376, -32'sd1667432, -32'sd1104333, -32'sd260646, -32'sd3833893, 
    -32'sd2939036, -32'sd2235985, -32'sd420899, -32'sd2286327, 32'sd183443, -32'sd976891, 32'sd1612842, -32'sd3545687, 
    -32'sd554416, 32'sd3919660, -32'sd48306, -32'sd1362209, 32'sd3937738, 32'sd1400424, -32'sd846154, 32'sd1976782
    };
    task set_inp_1;
        input integer task_int_len;
        input integer task_int_inv_len;
        begin
            for (n = 0; n < task_int_inv_len; n = n + 1)
                for (m = 0; m < task_int_len; m = m + 1) begin
                    temp_inp[((((n*2)*task_int_len)+m)*32)+:32] <=
                        temp_inp[((((n*2)*task_int_len)+m)*32)+:32] +
                        temp_inp[((((n*2)*task_int_len)+task_int_len+m)*32)+:32];
                    temp_i1[(((n*task_int_len)+m)*32)+:32] <=
                        -zetas[(((2*task_int_inv_len)-n-1)*32)+:32];
                    temp_i2[(((n*task_int_len)+m)*32)+:32] <=
                        temp_inp[((((n*2)*task_int_len)+m)*32)+:32] -
                        temp_inp[((((n*2)*task_int_len)+task_int_len+m)*32)+:32];
                end
        end
    endtask

    task set_inp_2;
        input integer task_int_counter;
        for (n = 0; n < 128; n = n + 1) begin
            temp_i1[(n*32)+:32] <= temp_inp[(((task_int_counter*128)+n)*32)+:32];
            temp_i2[(n*32)+:32] <= f;
        end
    endtask

    task set_out_1;
        input integer task_int_len;
        input integer task_int_inv_len;
        begin
            for (n = 0; n < task_int_inv_len; n = n + 1)
                for (m = 0; m < task_int_len; m = m + 1)
                    temp_inp[((((n*2)*task_int_len)+task_int_len+m)*32)+:32] <=
                        temp_o2[(((n*task_int_len)+m)*32)+:32];
        end
    endtask

    task set_out_2;
        input integer task_int_counter;
        for (n = 0; n < 128; n = n + 1)
            temp_inp[(((task_int_counter*128)+n)*32)+:32] <= temp_o2[(n*32)+:32];
    endtask

    genvar i;
    generate
        for (i = 0; i < 128; i = i + 1)
        begin: fqmul_32bit
            fqmul_32bit new_fqmul_32bit (
                .clock(clock),
                .reset(reset),
                .start(new_fqmul_32bit_start),
                .done(new_fqmul_32bit_done[i]),
                .a(temp_i1[(i*32)+:32]),
                .b(temp_i2[(i*32)+:32]),
                .reduce(temp_o1[(i*32)+:32])
            );
        end
    endgenerate

    assign new_fqmul_32bit_final_done = &new_fqmul_32bit_done;

    assign rd_ready = temp_rd_ready;
    assign rd_done  = temp_rd_done;
    assign done     = temp_done;
    assign wr_done  = temp_wr_done;
    assign out      = temp_out;

    always @(*) temp_o2 = temp_o1;

    // ======= FSM ch�nh =======
    always @(posedge clock)
        if (reset)
            state <= IDLE;
        else
            state <= next_state;

    always @(*) begin
        case (state)
            IDLE:        next_state = PRE_RD_INP;
            PRE_RD_INP:  next_state = start ? RD_INP : PRE_RD_INP;
            RD_INP:      next_state = CALC_1;
            CALC_1:      next_state = CALC_2;
            CALC_2:      next_state = new_fqmul_32bit_final_done ?
                                      ((len << 1) <= 9'd128 ? CALC_1 : CALC_3) : CALC_2;
            CALC_3:      next_state = CALC_4;
            CALC_4:      next_state = new_fqmul_32bit_final_done ?
                                      ((counter + 1'b1 < 2'd2) ? CALC_3 : WR_OUT) : CALC_4;
            WR_OUT:      next_state = DONE;
            DONE:        next_state = IDLE;
            default:     next_state = IDLE;
        endcase
    end
    always @(posedge clock) begin
        case (state)
            IDLE: begin
                counter <= 0;
                temp_rd_ready <= 0;
                temp_rd_done  <= 0;
                temp_done     <= 0;
                temp_wr_done  <= 0;
                temp_out      <= 0;
                len <= 9'd1;
            end
            PRE_RD_INP: begin
                if (start) temp_rd_ready <= 1;
            end
            RD_INP: begin
                temp_inp <= inp;
                temp_rd_ready <= 0;
                temp_rd_done  <= 1;
            end
            CALC_1: begin
                new_fqmul_32bit_start <= 1;
                case(len)
                    9'd1:   set_inp_1(1,128);
                    9'd2:   set_inp_1(2,64);
                    9'd4:   set_inp_1(4,32);
                    9'd8:   set_inp_1(8,16);
                    9'd16:  set_inp_1(16,8);
                    9'd32:  set_inp_1(32,4);
                    9'd64:  set_inp_1(64,2);
                    9'd128: set_inp_1(128,1);
                    default:set_inp_1(0,0);
                endcase
            end
            CALC_2: begin
                new_fqmul_32bit_start <= 0;
                if (new_fqmul_32bit_final_done) begin
                    case(len)
                        9'd1:   set_out_1(1,128);
                        9'd2:   set_out_1(2,64);
                        9'd4:   set_out_1(4,32);
                        9'd8:   set_out_1(8,16);
                        9'd16:  set_out_1(16,8);
                        9'd32:  set_out_1(32,4);
                        9'd64:  set_out_1(64,2);
                        9'd128: set_out_1(128,1);
                        default:set_out_1(0,0);
                    endcase
                    len <= len << 1;
                end
            end
            CALC_3: begin
                new_fqmul_32bit_start <= 1;
                case(counter)
                    2'd0: set_inp_2(0);
                    2'd1: set_inp_2(1);
                    default: set_inp_2(0);
                endcase
            end
            CALC_4: begin
                new_fqmul_32bit_start <= 0;
                if (new_fqmul_32bit_final_done) begin
                    case(counter)
                        2'd0: set_out_2(0);
                        2'd1: set_out_2(1);
                        default: set_out_2(0);
                    endcase
                    counter <= counter + 1'b1;
                end
            end
            WR_OUT: begin
                temp_out <= temp_inp;
                temp_done <= 1;
                temp_wr_done <= 1;
            end
            DONE: begin
                temp_done <= 0;
            end
            default: begin
                counter <= 0;
                new_fqmul_32bit_start <= 0;
                temp_inp <= 0;
                temp_i1 <= 0;
                temp_i2 <= 0;
                temp_rd_ready <= 0;
                temp_rd_done <= 0;
                temp_done <= 0;
                temp_wr_done <= 0;
                temp_out <= 0;
                len <= 9'd2;
            end
        endcase
    end
endmodule
