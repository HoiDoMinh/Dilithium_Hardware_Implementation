
module poly_pointwise_montgomery(
    input signed [8191:0] a_in,
    input signed [8191:0] b_in,
    output signed [8191:0]c_out
    );
    
    localparam N = 256;
    
    wire signed [31:0] a [0:N - 1];
    wire signed [31:0] b [0:N - 1];
    wire signed [31:0] c [0:N - 1];
    wire signed [63:0] mult64 [0:N - 1];
    
    generate
        genvar x;
        for (x = 0; x < N; x = x + 1) begin
		    assign a[x] = a_in[32 * x + 31:32 * x];
		    assign b[x] = b_in[32 * x + 31:32 * x];
		    assign mult64[x] = a[x] * b[x];
		    montgomery_reduce montgomery_reduce(.a(mult64[x]), .t(c[x]));
		    assign c_out[32 * x + 31:32 * x] = c[x]; 
		end
	endgenerate
    
endmodule