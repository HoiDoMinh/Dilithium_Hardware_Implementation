
`timescale 1ns/1ps
`include "byte_and_print.vh"

module tb_pack_sk;
    reg  [255:0]     rho_in;      // 32 bytes
    reg  [255:0]     key_in;      // 32 bytes
    reg  [511:0]     tr_in;       // 64 bytes (TRBYTES = 64)
    reg  [49151:0]   t0_in;     // 6 polys � 8192 bit
    reg  [40959:0]   s1_in;       // 5 polys � 8192 bit
    reg  [49151:0]   s2_in;       // 6 polys � 8192 bit
    wire [32255:0]   sk_out;   
    pack_sk dut(
    .rho_in(rho_in),      
    .key_in(key_in),     
    .tr_in(tr_in),      
    .t0_in(t0_in),       
    .s1_in(s1_in),      
    .s2_in(s2_in),      
    .sk_out (sk_out)      
    );


    wire [7:0] sk_bytes [0:4031];

    integer i;

    `BYTE_ASSIGN_GEN(SK, 4032, sk_out, sk_bytes)


    initial begin

        //
assign  rho_in = 256'h449e6340f762807b7675c26c548f69d84e7c623176dc341ee7bc8bc4b13f77e5;
assign  key_in = 256'he919c95dee122be585439e9350a9310e0308c433f9a12bac2e4227759ffd1195;
assign tr_in = 512'hea1d6a0dad5081a983e68f6d5e6abd327aed3f6c8cde5b7884a49f7e8c3397836440998a99bd820f3d51e471875fb94c6a180c3782615f2ae0ff97a9a1c28cd3;
assign t0_in = 49152'h00000b7300000f7000000c3200000ad3000004d900000ae000000220fffff9dffffffb30000000800000087900000efc00000487fffffa54fffff6c30000000bfffff7a9fffff5b40000042afffffc86fffffb93fffff8f8fffff7e800000ea80000088afffff496fffffc00fffff4da00000643ffffff1b00000a4300000ceafffff46600000e42fffff3f8fffff07cfffffa87fffffcaeffffff330000095b00000e13fffff785000008aa0000065500000dbd00000069fffffb6b00000132fffff68d000004d80000043dfffff6a5fffffa2d0000030afffffa8ffffffb5ffffff8a00000014d000005a6fffff650000004c7fffffd19000002b200000445fffffb33ffffff5800000f5afffffeb3000007f7fffffccfffffff3400000099fffff8390000096dfffffc41000003fafffff7a2fffff73dfffff686000006dffffffaac000007ddfffffea6fffff42500000a66000003d8fffff25bfffff880fffffca60000005a000004d2fffffe880000040900000fe9fffff750fffff182fffff2f2000006a90000030efffff5b800000a56fffff4d6fffff79100000262fffff1b1000004c8fffffc2dfffff782000002b0fffff13400000fa70000072700000ca20000053efffff6e60000037900000ef1000003ceffffff5e00000044fffff2e8fffffc7afffff762000009f0fffff505fffffed800000863fffff1fcffffff24000005aa000004dd000004bf0000005dfffff2e900000ce6fffff936fffff1fefffff149fffffd8bfffff9ddfffffdd2000009a500000ab6ffffffacfffff7c600000819fffff8c4fffffceefffff3c9fffff15efffff323fffffb54fffff7d3000001cdfffff20efffffa8efffff368fffffe05fffffa37fffff47dfffff15f00000e8400000eeefffffa2c00000edffffff2e100000f5cfffff57cfffff29afffffd5dfffff5910000032200000f2bfffff9e0000009cbfffff0e90000052efffff7c2fffff9ff00000d8800000c0e000008a8fffffb54000006b300000b95fffff58a0000026cfffffe200000090000000d6dfffff66cfffff63d00000abafffff2cb00000b0300000b5dfffffca400000e1a00000f8fffffffae000001bafffffa9bfffffde80000030500000023000001b6fffff57100000fc5ffffffad000003d3ffffff1800000fec00000950fffff10cfffff4520000079d00000b88fffff047000005c70000027c00000cea00000e8f00000dccfffff9b100000d54fffff1e100000f240000070600000dbc0000093a00000000000002f900000d8cffffff1800000d3d00000556fffffc3bfffff411000006cf000005120000031400000d0afffff345fffff92a00000f0600000fb3fffffa55fffffc7efffff46efffff5f3fffffa9300000a3200000646fffffee7000000cbfffff08000000fabfffff041fffff5c60000002500000671fffffc1100000e8300000fc70000094c00000ff4fffff3bdffffff2cffffffe5fffff429fffff733fffffa0e0000016afffffb950000099a0000038dfffffee500000ed200000af1fffff3a200000a8400000b4d0000071400000416fffffb4c00000a59fffff10300000a4500000ea60000008c00000623000005f6fffff35cfffff978fffff002000001a9fffff022000009f1fffff032000006a2fffff4670000070dfffff0fffffff34efffff2b300000930fffff63dfffffe68fffff211000001e6fffff0bcfffff815fffff804fffff5af0000099800000795fffff83400000f9100000849fffff3f200000dfb000009e8fffff059fffff30afffffb6e000002cefffff791000007fc00000148fffff1e800000f4cffffff3bfffff2da000009d5fffff283fffff7560000002f00000464fffffd810000000cfffff58300000381ffffffdefffff1e300000918000006a4ffffffe9000009d7000004bffffff8e2fffffaebfffff47100000243000002c60000062500000b340000024700000a300000089efffff309000009f800000f7cfffff1db00000a32fffff920fffffa32000008c7fffffc5e000005c300000f47fffff4ae00000df20000033200000b3c00000bbb00000ba7fffff296000006ef00000e29fffff747fffff413fffffa38fffffec300000b08000008bb00000030fffff2c0fffff65cfffff56600000527fffff491fffffd66fffffdcf00000a700000064c000006dc0000050f00000ac80000048dfffff57f000009470000071d00000f1bfffff080ffffffc7000007ee000003fc000003a8000008dffffff21a00000247000004cb000000fcfffff441fffffa240000085500000d150000092cfffff8f0fffff7b1fffff07200000b45fffff04bfffff5e2fffff569fffffe62ffffff52fffff7da00000662fffffba400000cf600000d6400000218fffff0e700000bfffffff6d9ffffff20000001fffffff6ca000004a2000004ab000002a2fffff753fffff685fffff66b000006dc00000cb2ffffffe6fffff0e0000002cb00000be9fffff8ac00000081000007d5000003f400000b7b00000631fffff325fffff613000001f6fffff88100000c72fffff998000009b3fffff6e3000008eafffffbc5ffffffcf00000318fffffa700000028efffffe27fffff852ffffff12fffff19a00000cd0fffff10200000882000007790000061000000856fffff756000003c9fffffcbe00000aa5000000e6fffff1a60000024cfffff209fffff17b00000b770000017a0000091c000006f600000428fffff7bdfffffd520000099d00000b3e0000028a0000070f00000a9efffff493fffff198000006acfffff30ffffff47dfffff99bffffffcffffffa9e000000d4fffff2a7000009d2fffff8bcfffff3ad0000050d000002ca0000023bfffff67cfffff155fffff0e90000038cfffff690fffff0420000032d0000063b000008bd000007effffffa390000090f0000097400000cf6fffff17c00000ef700000a74fffff820000006a900000c8d00000af6fffff96800000362fffff7f400000290000002cefffff582fffff1c800000314fffffe2cfffff3290000057afffffdc1000006e6fffffb20fffff51cffffff9d00000d8dfffffbbcfffff1e9fffff79afffffe40fffffb8a0000078efffff46dfffff02ffffffbfefffff92e000009a0000004a7fffffdfffffff63a00000e96fffff24200000ef4fffffcc2fffffa690000093afffffc2dfffff453000003af000002e10000026d00000711fffff517fffff47a00000c1400000e54fffff5de00000222000007410000082bfffff54cfffff03300000cb60000076700000b79fffffc7ffffff6d0fffff278000002da00000319fffff4f50000002dfffff113fffffda1fffff18100000296fffff3a3fffffd0ffffff69a00000a0000000889fffff3ccfffffb82fffff66afffff1b9ffffffa6fffff63dfffff072ffffff4900000a3e00000f82fffffc32fffff18e000002a200000926000008fcfffffa870000083f000001c2000002d3fffffb7efffffc2afffff15ffffffb6afffff9e700000506fffff6d600000696fffff815fffffb0afffffb65fffff20700000d47fffff98b0000093700000a83fffff45afffff20700000b470000021600000d5a00000fdb000005d8fffffa4f000001bffffff7c9fffff7b8fffff100fffffd5b000008430000053bfffff3ec00000ec0000001d8fffffd56fffff4e4fffff9460000036900000bc4fffff6440000064b000009d5000009b4fffff3b00000060800000771fffff99d00000f29000007a8fffff1edfffff00efffffbb6fffff5e900000afcfffffde5ffffff3bfffff94efffffe02fffffd6cfffff774ffffff44fffffebf000000db0000070efffffc1efffff7b1fffff2acfffffaaafffffcd60000099b000005b600000fd6fffff46800000d71fffff38f00000e7600000eecfffffb7f00000cf20000056afffffcdcfffffe3d00000cd10000019cfffff30700000d8900000678fffff7f6000005b0fffffa89fffff654fffffdd50000079f00000c72fffff4c3000009b100000a07fffff394fffffceffffff403fffff85afffffa76fffff9a700000106fffff5a0fffff2e50000028c000006b4000002f3000008f9fffffa19000002affffff62dfffff9cffffff0b0000005e600000cf600000b34fffff70d00000534fffff4bdfffff705fffff04bfffff3c6fffff813fffff347000009e9fffff448fffffe10fffff2d000000491fffffb8bfffff9cdfffff68b0000095cfffff96ffffff53b0000070d00000fdafffff84cfffff7c5000006f3000000f80000047b00000457fffff0e700000c8b00000cb5fffffca8fffffaf6fffffedafffff82dfffffc6a000002970000048a000007ba00000175fffffa420000003efffffe5cfffff48afffffc64fffff52d00000366000000d2000008c0ffffff6a0000024800000b90fffffdbf00000ee50000037300000465fffff76a00000731fffff0f3fffffc7bfffffb2100000290fffff3580000009800000c920000099cfffffe7dffffff19fffffb2afffff4890000042f000003b400000e69fffff08b000008050000099cfffffa81ffffff1d000003e600000ee9fffff0bffffff07500000bbdfffff274000004dbfffff79efffffd1ffffff02d00000aeafffff47400000a79fffff3b7000000e10000053800000bb70000030600000af900000ef7fffff606000002a1fffff51b000000fefffff4e1fffffef60000044600000db500000d1dfffffdbd00000b970000047a00000b3efffff1c3fffff1ee000004e000000571000007d500000b42fffffa74fffffa84fffffdecfffff13800000578000003c0fffffbc3fffff7a3000002fd000002050000060400000d2d0000053cffffffdefffff01cfffff4b500000f22fffffee2ffffff6900000039fffff4c1000008d200000113fffff85400000a5efffff31100000805000009b200000d31fffff4aefffff71200000119fffff96efffff6f600000ad2ffffff38fffff6b2fffff8540000003cfffffa95fffff6e4fffff2070000085d00000c46fffff6d8fffffe47fffff033000005750000016600000706fffff0c100000cdd0000090200000311fffff56400000f91000000d800000066fffffacffffffe43ffffff09fffff3effffffe17fffff451fffff49b0000089b0000026700000e64fffff2d2fffff653000006f9fffff04b00000b3cfffff8e60000006a0000084b00000ed500000b18ffffffbe00000e080000092dfffffc8f000000c5fffffa8f0000017e0000068b00000b3000000510000004f50000032200000040fffffe9200000cec00000154fffff25400000b8dfffffc9c0000038300000bc9fffff590fffffcac00000709fffff17c00000718fffff74dfffffdccfffff4a700000100fffff4be00000393fffff8f8fffff9f0fffffdca00000847fffff59d00000e0500000713000007a1fffff1ac0000075500000f8100000f24fffffabefffff146fffff7dafffffb9effffff55fffffee2fffffec9fffff5b8fffffb87fffffacefffffe52fffff89ffffff361fffffafcfffffe7d000003fbfffff439fffffdcbfffffd9efffffdc9fffff8a2fffffb2f00000631fffff458fffffb31fffff79400000e75fffffb0a00000438fffffc820000067000000d9f000009edfffff60700000e050000066500000670000008a0000007d2fffff73ffffff1280000063900000da50000007d00000463000009ddfffffed900000cdcfffff50bfffff9d5000003920000029100000eaefffffecf00000f3200000ddafffff3cb000007f400000953fffffbc8fffffcfbfffff040fffffa1b0000072800000b83ffffff96fffffa55fffffcedfffff7db000006f9000001a9000006e4fffff923fffffc0c00000abf0000031f000009dfffffff2ffffffa33000001880000008efffffa7f00000330fffff3bb00000c79fffff8b6fffff56900000f6dfffff14afffff4fefffffb01fffff7f0fffff907fffff7cffffff61900000376fffffc0bfffff997fffff049fffffa1f000002c6000005a8fffff663fffffb970000090efffffc84fffff53000000537000005d30000086900000af700000ba80000079400000654fffffe2b00000126fffff9a2ffffff4afffffae9fffff18d00000cea00000eb5fffffc57fffffd0ffffffd98ffffff5a0000065ffffff994fffffda1fffffad0fffff926000009bc00000385ffffffbafffff59dffffff1bfffffa320000070a00000d3bfffffd2ffffff1fc00000672fffffc80fffff69afffff50efffff1490000047bfffffd4bfffff81e000003b8fffff0d1fffff530000003adfffffc7dfffffe77000008080000050d00000c58000004fe00000828fffffcb4fffff3b6000005a60000004cfffff7d3fffff22cfffff78b00000fa7fffff37800000319fffff8c9000008e200000f64fffff4ec000004d000000439fffff82ffffffc6efffff622fffff3fa00000876fffff896fffff8e5000003a7fffff471fffffd6affffffbffffffdc60000014cfffff26e000004ff00000c69fffff266fffff8250000024600000412fffffee800000d74fffff47700000e1dfffff85000000cd500000d83fffffa4100000219000008b8fffff7d100000becfffff2460000005a000000f5fffff7a8fffffbaf00000e5000000bd4fffffbf0fffff213fffffe6800000aecfffffb1f000005a700000c89fffff26100000f73fffff4d5fffffd67fffff5c500000b10fffff19ffffff00a000003d5ffffff21000009e700000c4cfffffb6f00000d84fffff96800000618fffff3c8000000f4ffffffacfffffb000000080c00000721ffffff97fffff6160000049c00000d2e00000ba2ffffffc8fffffde5fffff422fffffa28fffffe69fffff6d0fffff3cbfffff09dfffffd5b00000a60fffff2ee0000076f00000eb600000069fffff493000002a9000003c4fffff394000007a30000055600000c8dfffff98200000b98fffff72ffffffc0900000ac7fffff749fffff345fffff6ac00000c170000048bfffff45cffffffd6fffff7f900000618000001e0000001e3fffffacb0000016ffffffb2b000000290000090afffffd45fffff345fffff1fffffff57a000000b900000cccfffffa0600000743000002c3fffff5e6fffffd500000072700000dd600000d7cfffff478000005290000008100000a03ffffffc300000a50fffffadefffff61f00000e1effffff54000005ac0000063ffffffb4ffffff88500000a0f00000f7600000c85fffffc21fffffcfcfffffac0fffffc0b00000b2efffff17c00000a4effffff3a00000f31fffffd0afffffd52fffffbdbfffffbb2fffffb3300000f8200000864fffffeda00000212fffff00100000add00000acafffffcf200000beafffff77b0000043300000ee5fffff14400000dbbfffffb75000009b4fffffcf9fffff5b1fffff7bdfffff744fffff94500000f1cfffffcc200000706000002ae0000057700000512fffff895000008b2000000a300000f9e0000096e0000088a000001f9000007c5fffff5e500000b7efffff69a0000099a00000d9200000267fffffe53fffff5de00000d95fffffca1fffff317fffffea400000a01fffff29900000372fffff924fffff24f0000068c00000a8d000000e600000359fffffad3fffffa900000078300000d69fffff4df0000090c0000039100000e67ffffff85fffff0f8fffff59c00000a26000000ba0000075c00000313fffff2fa0000063600000ccafffff87dfffff63dfffffdcafffff206fffffb54fffff5e9fffffb6f0000000afffff64c0000076600000d37fffffd42fffffb0afffffc8b0000055f00000a23fffff0b800000dc3fffffd0b000006fefffff59e0000091affffff1bfffffe58fffff5fafffffe9c00000a77fffffc5c0000039d000000270000062a000009fefffff2310000057200000447fffffd93fffff1ce000004eb00000dec000001c80000014c000007d5000008dd000003fffffff57700000b35000009fe000005cbfffff0affffff37900000398fffff11ffffff3cafffffd87fffff6c8fffff3b700000f2cffffff0d000001ddfffff16900000bb9fffffdfffffff7e400000db1fffff0f00000006100000a2e00000c38000008f7fffff37b00000e27000008bdfffff1ba0000011bfffffc8e000006c300000185fffff2cdfffff7b200000fb800000e6dfffffe11fffff52900000233000006b7fffffb19fffff8770000066c00000983fffff1dc00000526fffffbabffffff5dfffff15afffffa6f000003ccfffff5c6000008d0ffffface000003850000033ffffffe8b00000ed7000006f50000098900000e56000006c4fffff15e00000c5500000cb9fffff6ac00000b4400000d11fffffabd0000012cfffff36b00000f7cfffffe100000071e000005830000084a00000b5a000006f5000007860000045afffff8bcfffffbaffffff83100000e18fffffe98000008dd00000648fffff383fffff3b600000e3300000f830000027f000005cbfffff185000000b4;
assign s1_in = 40960'h0000000000000001ffffffff0000000100000001fffffffc000000000000000200000000fffffffe0000000100000001fffffffd000000000000000300000000fffffffdfffffffdffffffff00000002fffffffc000000000000000100000000000000040000000000000004fffffffc00000004ffffffff00000003fffffffcfffffffc0000000000000002fffffffd000000040000000100000003fffffffdfffffffe00000002000000010000000400000000fffffffe00000003fffffffdffffffff0000000400000002fffffffdfffffffe00000001fffffffcfffffffcfffffffe000000000000000000000002fffffffdfffffffd000000040000000000000003fffffffdfffffffefffffffcfffffffe0000000000000003000000010000000400000001fffffffdfffffffffffffffc00000000fffffffffffffffe00000003fffffffffffffffe00000004fffffffd00000003fffffffefffffffcfffffffd000000020000000000000001fffffffc0000000400000004fffffffcfffffffffffffffefffffffd00000003000000020000000000000004fffffffefffffffffffffffc00000004fffffffe000000040000000400000000fffffffc000000020000000200000003fffffffe0000000400000004fffffffd0000000400000001ffffffff00000003fffffffd00000002000000030000000300000004000000030000000200000001fffffffc000000000000000000000000fffffffe0000000300000001fffffffffffffffcffffffff0000000400000001fffffffdfffffffe0000000000000002000000030000000300000002fffffffc0000000300000001000000010000000400000001000000030000000200000004fffffffe0000000000000000ffffffff00000002ffffffff00000003fffffffc00000003fffffffe0000000200000004fffffffffffffffd000000000000000200000001fffffffe00000003fffffffefffffffffffffffdffffffff00000003fffffffd000000000000000400000003fffffffdfffffffffffffffc000000020000000200000001fffffffffffffffd00000003fffffffcfffffffffffffffeffffffff00000000ffffffff00000002fffffffdffffffff000000030000000200000004fffffffe00000003000000030000000200000000fffffffdfffffffe0000000000000004ffffffff00000004fffffffffffffffffffffffdfffffffffffffffcfffffffd0000000400000004ffffffff000000020000000400000000fffffffc00000002fffffffdffffffffffffffff00000003fffffffd000000000000000300000000fffffffc000000040000000400000004fffffffffffffffc00000001fffffffe00000002fffffffcfffffffeffffffff0000000300000000ffffffff0000000100000002ffffffff00000000fffffffdfffffffffffffffcffffffff00000004fffffffdfffffffc0000000000000002fffffffefffffffc00000002fffffffe000000010000000000000004fffffffd00000002fffffffefffffffffffffffcfffffffdfffffffdffffffff00000000fffffffefffffffd00000000ffffffff000000040000000100000000fffffffdfffffffe000000000000000100000004000000020000000400000002ffffffffffffffff00000001fffffffd0000000300000002fffffffd0000000200000003fffffffe00000003fffffffc0000000200000000000000040000000100000002fffffffdfffffffd00000004fffffffcfffffffffffffffc00000004ffffffff00000002fffffffeffffffff0000000100000001fffffffe00000000fffffffc00000004fffffffefffffffffffffffffffffffefffffffe00000001fffffffd00000000ffffffff00000003fffffffffffffffcfffffffe0000000200000003fffffffe0000000300000000000000040000000000000003fffffffefffffffc000000040000000400000000fffffffeffffffff00000002fffffffdfffffffefffffffe00000003000000010000000100000000fffffffcfffffffd0000000200000003fffffffffffffffdfffffffffffffffffffffffffffffffe0000000000000001fffffffffffffffffffffffd00000000fffffffffffffffcfffffffc00000002fffffffe00000001fffffffdfffffffe0000000000000002fffffffdfffffffcfffffffe00000001fffffffe00000000fffffffffffffffc00000001fffffffc00000003fffffffcffffffff00000003fffffffe0000000300000001fffffffd00000000fffffffefffffffc00000002ffffffff00000004ffffffff00000003ffffffff00000003fffffffefffffffffffffffcfffffffc00000002000000040000000200000001000000000000000100000000fffffffcfffffffd00000003fffffffdfffffffffffffffdfffffffd0000000200000003fffffffd00000001ffffffff0000000400000004fffffffffffffffd0000000400000002000000040000000000000002fffffffe00000003fffffffcfffffffc00000004000000010000000300000002fffffffffffffffe00000003fffffffc00000004fffffffc0000000200000002fffffffdffffffff00000003000000000000000300000002fffffffefffffffffffffffdfffffffefffffffc0000000400000002fffffffc0000000000000004fffffffe00000004fffffffe0000000400000004fffffffd00000000fffffffd00000002000000010000000000000004fffffffdfffffffcfffffffffffffffd00000003000000020000000000000000fffffffe00000003fffffffcfffffffcfffffffd00000004fffffffc00000002fffffffc000000010000000300000000fffffffcfffffffdfffffffd0000000100000003fffffffd00000001000000010000000200000004ffffffff00000004ffffffff0000000000000000fffffffdffffffff0000000200000004fffffffefffffffc00000003fffffffd000000000000000200000001fffffffd000000020000000100000000fffffffefffffffcffffffff00000003fffffffcfffffffd00000001fffffffd0000000100000002000000030000000200000000fffffffe0000000100000000fffffffd00000003ffffffff0000000100000002fffffffffffffffcfffffffdfffffffd00000003fffffffe0000000200000001ffffffff00000000fffffffefffffffefffffffffffffffdfffffffd000000010000000000000004fffffffe00000003fffffffd00000002fffffffefffffffeffffffff00000001fffffffcffffffff0000000200000002fffffffc0000000300000002fffffffefffffffd00000001ffffffffffffffff00000003fffffffc00000004fffffffd00000001ffffffff00000003fffffffcfffffffcffffffff0000000000000003fffffffc00000002fffffffcfffffffdfffffffefffffffffffffffffffffffefffffffffffffffeffffffff00000002fffffffdfffffffd0000000000000002fffffffd00000002fffffffe00000001fffffffc00000001fffffffdffffffff0000000100000003000000000000000100000000fffffffd0000000300000003fffffffefffffffe0000000100000002fffffffffffffffffffffffdfffffffc0000000200000000fffffffefffffffdfffffffefffffffe00000004fffffffdfffffffc0000000200000000fffffffcfffffffcfffffffd00000004fffffffefffffffdfffffffc0000000100000004fffffffcfffffffcfffffffefffffffd000000030000000300000004fffffffc00000002fffffffffffffffe0000000000000000ffffffff000000040000000200000001fffffffe00000002fffffffdfffffffdffffffff00000000fffffffd00000004fffffffc00000000fffffffefffffffc0000000400000001ffffffffffffffff000000030000000100000003fffffffefffffffd0000000400000002fffffffefffffffdfffffffcfffffffffffffffc0000000400000003fffffffd00000000fffffffcfffffffefffffffe000000000000000300000003ffffffff00000002fffffffffffffffd0000000100000002fffffffdfffffffe00000001fffffffefffffffeffffffff0000000000000002fffffffe000000000000000400000001fffffffcfffffffffffffffdfffffffefffffffefffffffdfffffffcfffffffdfffffffcfffffffdfffffffe000000040000000400000002fffffffdfffffffe0000000000000004fffffffcfffffffffffffffc000000040000000000000002fffffffd00000004fffffffd00000004fffffffefffffffe000000000000000300000000fffffffe00000001000000030000000100000003fffffffc0000000000000001fffffffe00000001ffffffff00000003fffffffd00000000fffffffffffffffeffffffff00000004fffffffc0000000000000004fffffffffffffffdfffffffc00000001fffffffefffffffffffffffe00000003fffffffefffffffffffffffefffffffe0000000000000002fffffffe00000003fffffffffffffffdfffffffffffffffd0000000400000000ffffffff0000000100000000fffffffcfffffffdfffffffd0000000300000002ffffffffffffffff00000002000000010000000000000003ffffffff0000000300000002000000000000000000000002fffffffe0000000200000000ffffffff00000001fffffffcfffffffd0000000200000004fffffffdffffffff0000000200000000fffffffe0000000100000002fffffffdfffffffcffffffff00000002fffffffc00000002ffffffff00000001fffffffcfffffffe0000000300000004fffffffdfffffffc00000001fffffffd00000000fffffffe00000000fffffffffffffffd0000000400000003000000040000000400000000fffffffc000000010000000300000001fffffffefffffffe00000004000000040000000400000001fffffffefffffffd000000020000000400000004fffffffd0000000100000004fffffffdfffffffc000000020000000100000003fffffffffffffffffffffffffffffffe0000000200000004fffffffe0000000100000001fffffffdfffffffc0000000100000002fffffffc0000000300000002fffffffeffffffffffffffff000000030000000400000001000000020000000100000001ffffffff000000040000000300000004000000030000000400000004fffffffcfffffffd0000000000000004fffffffd000000010000000200000002fffffffc0000000000000003fffffffffffffffffffffffcfffffffd000000040000000400000004fffffffc00000002fffffffffffffffffffffffcfffffffe0000000100000002fffffffd0000000300000003fffffffcfffffffd0000000000000001fffffffdfffffffc0000000200000002fffffffefffffffffffffffffffffffe00000000fffffffcfffffffc0000000000000004fffffffdfffffffefffffffc00000004000000000000000200000000fffffffffffffffe00000003fffffffefffffffdfffffffcfffffffcfffffffefffffffdfffffffcffffffffffffffff00000002fffffffd00000003fffffffd00000002fffffffffffffffdfffffffe00000004000000010000000300000002fffffffdffffffff00000002fffffffefffffffdfffffffd000000010000000300000003fffffffd00000000ffffffff00000000fffffffffffffffefffffffffffffffcffffffff0000000200000003ffffffff0000000000000001fffffffffffffffffffffffd00000004000000000000000200000001ffffffff00000000000000010000000200000002000000010000000300000002fffffffffffffffdfffffffffffffffd0000000000000004fffffffd0000000400000004ffffffff00000003fffffffffffffffc00000001fffffffcffffffff00000003fffffffc0000000100000001fffffffdfffffffd0000000400000000fffffffeffffffff00000004ffffffff00000002fffffffefffffffe000000010000000200000001fffffffdfffffffd00000003fffffffcfffffffffffffffdfffffffc00000002fffffffc00000001fffffffc00000000fffffffefffffffefffffffe0000000300000002fffffffefffffffd00000003fffffffffffffffffffffffc0000000300000003000000020000000300000001fffffffc00000004fffffffcfffffffd00000002fffffffc00000002fffffffefffffffe00000003fffffffcfffffffefffffffcfffffffdfffffffd00000001fffffffd00000002fffffffcfffffffe000000000000000400000001fffffffc000000030000000200000004fffffffeffffffff00000001fffffffe00000001000000010000000400000002000000020000000200000003fffffffdfffffffeffffffffffffffff000000010000000100000001fffffffd0000000400000000fffffffeffffffff00000000000000030000000000000003ffffffff000000010000000200000004000000000000000100000001fffffffd00000000fffffffcfffffffc0000000300000003fffffffc00000001fffffffffffffffe00000002fffffffffffffffc000000030000000400000002fffffffcffffffff0000000300000002fffffffcfffffffd00000003fffffffe000000040000000200000002fffffffdfffffffd00000004fffffffefffffffd00000000fffffffffffffffefffffffdfffffffe0000000000000001000000040000000000000002fffffffe000000040000000300000001000000030000000000000002000000010000000100000001fffffffcfffffffe00000002fffffffefffffffe00000004ffffffff0000000100000003fffffffc000000010000000000000004fffffffe00000000fffffffd000000030000000200000001ffffffff000000020000000000000000ffffffff00000002fffffffd00000000fffffffdfffffffffffffffcfffffffc00000004fffffffcfffffffdffffffff0000000100000002fffffffe000000030000000300000003fffffffe00000003;
assign s2_in = 49152'hfffffffffffffffcfffffffcfffffffc00000000fffffffd00000001000000020000000100000002fffffffefffffffefffffffd0000000200000001ffffffff0000000200000001fffffffe00000000fffffffcfffffffd00000002fffffffe00000004ffffffff00000001fffffffe00000003ffffffff00000003fffffffe000000040000000300000003fffffffcfffffffc000000020000000100000001fffffffe00000000fffffffffffffffe0000000100000001fffffffc0000000300000003fffffffe000000030000000200000003fffffffe00000002fffffffdfffffffe00000003000000010000000200000003ffffffff00000003fffffffcfffffffffffffffdfffffffe0000000300000002fffffffd0000000400000004fffffffcfffffffcfffffffe0000000100000004ffffffff00000003fffffffe0000000400000004000000020000000200000001ffffffff00000000fffffffc00000001fffffffd00000002fffffffd000000040000000200000004fffffffdffffffff000000010000000300000002fffffffdfffffffe00000004ffffffff00000000000000020000000400000000fffffffdfffffffc00000004fffffffdffffffff00000004fffffffe00000004ffffffff00000003fffffffdfffffffe0000000400000002fffffffc00000000ffffffff000000040000000000000001ffffffff00000004fffffffe00000000fffffffc00000000fffffffdffffffff0000000200000001ffffffff0000000000000004ffffffff00000002fffffffc00000004fffffffe00000004fffffffdfffffffd000000000000000100000003fffffffc0000000100000001fffffffc00000004fffffffefffffffefffffffffffffffd00000000fffffffeffffffff00000002fffffffe00000003000000030000000300000002ffffffff0000000200000000ffffffff00000002fffffffffffffffe000000030000000000000001fffffffffffffffe000000040000000200000001000000000000000100000000fffffffdfffffffe0000000200000003000000010000000300000003fffffffefffffffe00000001fffffffcfffffffcfffffffd000000020000000200000004fffffffffffffffefffffffd00000003fffffffc0000000400000003fffffffcfffffffc00000002fffffffd00000001ffffffff00000003000000040000000400000001fffffffe0000000300000003fffffffefffffffdffffffff00000004000000020000000000000003fffffffcffffffff0000000400000003000000020000000100000002fffffffdfffffffe0000000000000002fffffffdfffffffe00000003000000040000000000000001fffffffcfffffffffffffffd00000000fffffffcfffffffdfffffffe0000000300000002fffffffc000000020000000300000000000000020000000100000003fffffffd0000000000000004fffffffe00000000000000040000000000000000fffffffe00000002fffffffd00000001fffffffe0000000200000001ffffffff0000000000000002fffffffd00000002000000040000000400000002fffffffeffffffff0000000100000002fffffffd00000003fffffffd00000002000000010000000300000001fffffffe00000001fffffffefffffffdfffffffcfffffffefffffffffffffffd0000000100000001000000010000000200000000fffffffd00000003000000020000000000000002fffffffe0000000100000000fffffffc00000004fffffffffffffffc00000003fffffffe00000002fffffffdfffffffe00000003fffffffe0000000100000001fffffffc00000002fffffffefffffffe00000003fffffffe00000001fffffffd000000030000000400000002fffffffefffffffffffffffcfffffffe00000002000000030000000000000001fffffffc00000004fffffffdfffffffe00000000fffffffc00000000fffffffefffffffdfffffffe00000002fffffffd00000001fffffffe00000001fffffffc000000010000000200000001000000020000000000000000ffffffff000000020000000100000000000000020000000000000003000000000000000200000004ffffffff00000003000000020000000100000004fffffffe000000020000000200000004fffffffcfffffffc000000000000000200000000fffffffe0000000400000004fffffffcfffffffe00000002fffffffffffffffe00000004fffffffd00000003fffffffdfffffffd0000000400000001fffffffd000000020000000200000004fffffffd000000040000000200000000fffffffefffffffefffffffd00000000fffffffc000000010000000300000003fffffffc00000003000000010000000100000000fffffffdfffffffdfffffffefffffffefffffffe000000010000000100000003fffffffdfffffffe00000003fffffffc00000001ffffffff000000020000000000000001ffffffff0000000300000000fffffffeffffffff00000002fffffffefffffffd00000000fffffffffffffffdfffffffe00000002fffffffefffffffefffffffd0000000000000001ffffffff00000000fffffffe00000004fffffffc00000003000000030000000100000001fffffffe000000040000000400000003fffffffd0000000300000001fffffffc00000000000000030000000400000003fffffffdffffffff00000003fffffffffffffffc00000003fffffffffffffffd0000000100000000fffffffefffffffc0000000400000000000000020000000100000001ffffffff0000000000000004fffffffdfffffffc00000004fffffffe00000003ffffffff00000002fffffffefffffffc0000000100000003ffffffff00000003000000030000000100000003fffffffcfffffffefffffffe00000000fffffffc00000000fffffffefffffffe0000000400000002fffffffd00000000fffffffd000000010000000300000002fffffffcfffffffcfffffffc00000003fffffffcfffffffeffffffffffffffff00000004fffffffdfffffffc0000000200000002fffffffffffffffe00000004fffffffeffffffff000000010000000100000000fffffffd00000002000000040000000400000001fffffffffffffffc00000001000000010000000000000001fffffffcfffffffc00000003fffffffffffffffeffffffff0000000000000001fffffffd00000003fffffffffffffffcfffffffefffffffdfffffffd000000010000000100000004fffffffe00000003fffffffdfffffffd000000030000000100000003fffffffe00000004fffffffefffffffc000000000000000300000002fffffffcfffffffc00000002000000000000000100000002fffffffe0000000300000003fffffffd00000003fffffffc00000000fffffffffffffffefffffffc00000004fffffffc000000010000000200000000000000040000000000000000fffffffd0000000200000004fffffffeffffffff000000030000000100000001fffffffdffffffff000000030000000100000002fffffffcfffffffe0000000300000002ffffffff0000000000000001fffffffd0000000000000002fffffffc00000002fffffffcfffffffd000000030000000400000002ffffffff00000003fffffffefffffffe00000000fffffffffffffffefffffffe000000030000000300000003000000000000000000000000fffffffd00000002000000030000000300000000ffffffffffffffffffffffff0000000300000000fffffffffffffffe00000000fffffffd0000000200000003fffffffe0000000300000003fffffffcffffffff000000000000000300000000fffffffdffffffff000000020000000100000002fffffffe0000000400000002fffffffffffffffdfffffffeffffffff0000000100000003fffffffd00000002fffffffe00000000fffffffffffffffe00000003fffffffcffffffff0000000000000001ffffffff00000003fffffffffffffffc00000003fffffffdfffffffe0000000300000002000000030000000000000003fffffffefffffffc0000000400000000ffffffff00000003ffffffffffffffff0000000000000003000000000000000400000002fffffffc0000000000000002fffffffdfffffffdfffffffc0000000000000002000000020000000100000001fffffffcfffffffdfffffffdffffffffffffffff00000001fffffffcfffffffcfffffffffffffffdfffffffe0000000300000000fffffffdfffffffefffffffe000000040000000300000000fffffffefffffffe0000000400000003fffffffffffffffd0000000200000000fffffffd00000004fffffffdfffffffe0000000100000001fffffffd000000000000000000000003fffffffd00000003fffffffc00000001fffffffe00000000fffffffffffffffdfffffffe000000030000000200000002ffffffff00000002fffffffd00000004000000040000000400000004fffffffc00000004000000030000000000000000000000040000000100000002fffffffc00000004fffffffcfffffffeffffffff00000003fffffffdfffffffefffffffd00000003fffffffcffffffff00000000fffffffd00000000fffffffd000000030000000100000001fffffffc00000003fffffffd000000020000000400000002fffffffdfffffffc0000000000000000000000000000000200000004fffffffffffffffcfffffffc00000000000000010000000100000001fffffffd00000000fffffffeffffffff000000020000000100000000ffffffff00000001fffffffc00000001fffffffc00000000000000040000000100000002fffffffe00000001fffffffe00000001fffffffffffffffe0000000100000003fffffffeffffffff00000003fffffffcfffffffc0000000000000001fffffffe0000000300000003000000040000000200000001fffffffefffffffd00000002000000000000000100000000fffffffcfffffffcfffffffffffffffc00000003fffffffefffffffdfffffffd0000000000000003fffffffe00000004fffffffefffffffd00000004fffffffd00000001fffffffd0000000000000003000000030000000100000004000000020000000400000000fffffffdfffffffdfffffffe0000000300000001fffffffe000000000000000000000003fffffffffffffffc0000000100000002ffffffff0000000300000002000000000000000100000003ffffffff0000000100000000fffffffd00000001fffffffe0000000100000003fffffffcfffffffc00000001000000010000000000000002fffffffe00000001fffffffc0000000200000003ffffffff000000020000000100000004fffffffe00000003000000030000000100000004fffffffcfffffffc0000000300000002fffffffeffffffff0000000300000001fffffffe00000000fffffffefffffffcfffffffd00000003ffffffff0000000400000000fffffffe0000000000000000fffffffffffffffeffffffff00000000fffffffd0000000300000000fffffffd00000000000000010000000200000002fffffffc000000000000000300000001ffffffff0000000200000004fffffffe00000003fffffffc0000000400000000fffffffffffffffffffffffd00000004fffffffcfffffffc00000001fffffffc00000001fffffffc0000000200000002fffffffefffffffefffffffcfffffffe000000030000000200000004fffffffefffffffcfffffffcfffffffe00000000000000040000000200000002000000010000000300000001fffffffe0000000100000002fffffffefffffffd00000003000000010000000200000003000000000000000300000000000000040000000000000001fffffffe0000000200000003ffffffff00000002fffffffd0000000200000003ffffffffffffffff00000001000000010000000400000000fffffffd0000000300000000fffffffd00000002ffffffff00000002fffffffd00000001ffffffffffffffff000000000000000200000004ffffffff00000004fffffffcffffffff000000040000000300000000fffffffcfffffffffffffffcffffffff00000004fffffffd00000004fffffffeffffffffffffffff0000000200000000000000010000000100000002ffffffff00000001fffffffc00000000000000030000000000000001fffffffe00000002fffffffdfffffffeffffffff00000004fffffffe00000001fffffffefffffffe0000000300000003000000030000000000000002fffffffc00000001fffffffc000000030000000000000001000000010000000400000004ffffffff00000004fffffffc00000003fffffffe0000000200000000fffffffc00000004ffffffff0000000000000003fffffffefffffffc00000003000000020000000300000004fffffffdfffffffe0000000000000002000000030000000100000003fffffffc00000003fffffffc000000030000000400000003fffffffdffffffff00000000fffffffd0000000200000003fffffffe000000010000000000000000fffffffe0000000100000003fffffffc0000000300000004fffffffc0000000400000001fffffffe00000001fffffffc00000001fffffffefffffffcffffffff00000003fffffffffffffffefffffffdffffffff0000000300000003fffffffc00000002fffffffc00000002fffffffe00000004ffffffff00000004fffffffe0000000000000001ffffffff00000000fffffffe00000000000000030000000100000003fffffffcfffffffffffffffe00000003000000000000000300000002ffffffff000000010000000200000004fffffffffffffffd00000003fffffffdfffffffdfffffffd0000000300000001fffffffe0000000300000001fffffffc0000000400000003fffffffe00000004fffffffe00000000000000030000000400000001000000020000000200000003fffffffffffffffcfffffffc0000000300000000000000020000000100000004fffffffc0000000100000001ffffffff0000000000000002fffffffe0000000100000002fffffffe00000000fffffffd00000002000000000000000000000000fffffffefffffffc00000003fffffffd0000000100000001fffffffc00000001000000030000000400000001fffffffcfffffffdfffffffffffffffc00000001000000040000000100000004fffffffefffffffe00000001000000010000000300000000fffffffcfffffffeffffffff000000020000000000000004fffffffefffffffe0000000200000002fffffffdfffffffdfffffffd00000004fffffffd00000004fffffffcfffffffffffffffd00000004fffffffc0000000400000003fffffffdfffffffe0000000200000002fffffffcfffffffefffffffe0000000300000004fffffffe000000000000000200000000fffffffefffffffefffffffc00000002fffffffd00000001ffffffff000000030000000000000003fffffffc000000010000000000000003fffffffd0000000100000003fffffffc00000002fffffffe0000000200000004fffffffcffffffff000000000000000100000004fffffffefffffffdfffffffcfffffffc0000000200000002000000020000000400000003ffffffff00000003000000030000000400000004fffffffd00000001fffffffe00000001fffffffefffffffd00000003fffffffd00000003000000030000000100000001ffffffff00000002fffffffe0000000100000004fffffffefffffffd00000000fffffffc000000030000000400000001fffffffffffffffffffffffe00000001fffffffdfffffffdfffffffe0000000400000002fffffffcfffffffcfffffffd0000000200000004fffffffcfffffffcfffffffc00000001fffffffffffffffefffffffefffffffc0000000100000004000000010000000200000003fffffffefffffffeffffffff00000004000000010000000000000001ffffffff0000000200000002000000000000000400000003fffffffe00000000fffffffdffffffff00000002000000030000000100000001fffffffdffffffff00000004fffffffffffffffffffffffe00000003fffffffc00000004fffffffcfffffffc00000003fffffffcfffffffd00000001fffffffe00000002000000010000000200000004fffffffd00000000fffffffe00000002000000010000000300000002fffffffeffffffff0000000300000000fffffffd00000002000000010000000000000004fffffffe00000003ffffffff00000001fffffffd000000040000000300000004fffffffc0000000300000000fffffffffffffffe00000000fffffffc0000000100000000fffffffffffffffd0000000000000003fffffffefffffffcfffffffd000000030000000200000003fffffffd0000000100000001fffffffe0000000100000001000000010000000000000002ffffffff00000001;

        #10;

        `PRINT_HEX_ARRAY("sk_out (Verilog)", sk_bytes, 4032)

        $finish;
    end

endmodule